Simple Test Circuit
* Basic resistor divider for testing

V1 in 0 DC 5
R1 in out 1k
R2 out 0 1k

.op
.control
run
print all
.endc
.end
